`timescale 1ns/1ps

package tb_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import ahb_types_pkg::*;
  import ahb_uvm_pkg::*;

  // Tests
  `include "tb_tests.svh"
endpackage

